module Register8CE (input [7:0] I, output [7:0] O, input  CLK, input  CE);
wire  inst0_Q;
wire  inst1_Q;
wire  inst2_Q;
wire  inst3_Q;
wire  inst4_Q;
wire  inst5_Q;
wire  inst6_Q;
wire  inst7_Q;
SB_DFFE inst0 (.C(CLK), .E(CE), .D(I[0]), .Q(inst0_Q));
SB_DFFE inst1 (.C(CLK), .E(CE), .D(I[1]), .Q(inst1_Q));
SB_DFFE inst2 (.C(CLK), .E(CE), .D(I[2]), .Q(inst2_Q));
SB_DFFE inst3 (.C(CLK), .E(CE), .D(I[3]), .Q(inst3_Q));
SB_DFFE inst4 (.C(CLK), .E(CE), .D(I[4]), .Q(inst4_Q));
SB_DFFE inst5 (.C(CLK), .E(CE), .D(I[5]), .Q(inst5_Q));
SB_DFFE inst6 (.C(CLK), .E(CE), .D(I[6]), .Q(inst6_Q));
SB_DFFE inst7 (.C(CLK), .E(CE), .D(I[7]), .Q(inst7_Q));
assign O = {inst7_Q,inst6_Q,inst5_Q,inst4_Q,inst3_Q,inst2_Q,inst1_Q,inst0_Q};
endmodule

module Add8 (input [7:0] I0, input [7:0] I1, output [7:0] O, output  COUT);
wire  inst0_O;
wire  inst1_CO;
wire  inst2_O;
wire  inst3_CO;
wire  inst4_O;
wire  inst5_CO;
wire  inst6_O;
wire  inst7_CO;
wire  inst8_O;
wire  inst9_CO;
wire  inst10_O;
wire  inst11_CO;
wire  inst12_O;
wire  inst13_CO;
wire  inst14_O;
wire  inst15_CO;
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst0 (.I0(1'b0), .I1(I0[0]), .I2(I1[0]), .I3(1'b0), .O(inst0_O));
SB_CARRY inst1 (.I0(I0[0]), .I1(I1[0]), .CI(1'b0), .CO(inst1_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst2 (.I0(1'b0), .I1(I0[1]), .I2(I1[1]), .I3(inst1_CO), .O(inst2_O));
SB_CARRY inst3 (.I0(I0[1]), .I1(I1[1]), .CI(inst1_CO), .CO(inst3_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst4 (.I0(1'b0), .I1(I0[2]), .I2(I1[2]), .I3(inst3_CO), .O(inst4_O));
SB_CARRY inst5 (.I0(I0[2]), .I1(I1[2]), .CI(inst3_CO), .CO(inst5_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst6 (.I0(1'b0), .I1(I0[3]), .I2(I1[3]), .I3(inst5_CO), .O(inst6_O));
SB_CARRY inst7 (.I0(I0[3]), .I1(I1[3]), .CI(inst5_CO), .CO(inst7_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst8 (.I0(1'b0), .I1(I0[4]), .I2(I1[4]), .I3(inst7_CO), .O(inst8_O));
SB_CARRY inst9 (.I0(I0[4]), .I1(I1[4]), .CI(inst7_CO), .CO(inst9_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst10 (.I0(1'b0), .I1(I0[5]), .I2(I1[5]), .I3(inst9_CO), .O(inst10_O));
SB_CARRY inst11 (.I0(I0[5]), .I1(I1[5]), .CI(inst9_CO), .CO(inst11_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst12 (.I0(1'b0), .I1(I0[6]), .I2(I1[6]), .I3(inst11_CO), .O(inst12_O));
SB_CARRY inst13 (.I0(I0[6]), .I1(I1[6]), .CI(inst11_CO), .CO(inst13_CO));
SB_LUT4 #(.LUT_INIT(16'hC33C)) inst14 (.I0(1'b0), .I1(I0[7]), .I2(I1[7]), .I3(inst13_CO), .O(inst14_O));
SB_CARRY inst15 (.I0(I0[7]), .I1(I1[7]), .CI(inst13_CO), .CO(inst15_CO));
assign O = {inst14_O,inst12_O,inst10_O,inst8_O,inst6_O,inst4_O,inst2_O,inst0_O};
assign COUT = inst15_CO;
endmodule

module Mux2x8 (input [7:0] I0, input [7:0] I1, input  S, output [7:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(S), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(S), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(S), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(S), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst4 (.I0(I0[4]), .I1(I1[4]), .I2(S), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst5 (.I0(I0[5]), .I1(I1[5]), .I2(S), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst6 (.I0(I0[6]), .I1(I1[6]), .I2(S), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'hCACA)) inst7 (.I0(I0[7]), .I1(I1[7]), .I2(S), .I3(1'b0), .O(inst7_O));
assign O = {inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module Decoder4 (input [3:0] I, output [15:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
SB_LUT4 #(.LUT_INIT(16'h0001)) inst0 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h0002)) inst1 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h0004)) inst2 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h0008)) inst3 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h0010)) inst4 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h0020)) inst5 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h0040)) inst6 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h0080)) inst7 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst7_O));
SB_LUT4 #(.LUT_INIT(16'h0100)) inst8 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst8_O));
SB_LUT4 #(.LUT_INIT(16'h0200)) inst9 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst9_O));
SB_LUT4 #(.LUT_INIT(16'h0400)) inst10 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst10_O));
SB_LUT4 #(.LUT_INIT(16'h0800)) inst11 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst11_O));
SB_LUT4 #(.LUT_INIT(16'h1000)) inst12 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst12_O));
SB_LUT4 #(.LUT_INIT(16'h2000)) inst13 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst13_O));
SB_LUT4 #(.LUT_INIT(16'h4000)) inst14 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst14_O));
SB_LUT4 #(.LUT_INIT(16'h8000)) inst15 (.I0(I[0]), .I1(I[1]), .I2(I[2]), .I3(I[3]), .O(inst15_O));
assign O = {inst15_O,inst14_O,inst13_O,inst12_O,inst11_O,inst10_O,inst9_O,inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module And2x16 (input [15:0] I0, input [15:0] I1, output [15:0] O);
wire  inst0_O;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_O;
wire  inst9_O;
wire  inst10_O;
wire  inst11_O;
wire  inst12_O;
wire  inst13_O;
wire  inst14_O;
wire  inst15_O;
SB_LUT4 #(.LUT_INIT(16'h8888)) inst0 (.I0(I0[0]), .I1(I1[0]), .I2(1'b0), .I3(1'b0), .O(inst0_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst1 (.I0(I0[1]), .I1(I1[1]), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst2 (.I0(I0[2]), .I1(I1[2]), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst3 (.I0(I0[3]), .I1(I1[3]), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst4 (.I0(I0[4]), .I1(I1[4]), .I2(1'b0), .I3(1'b0), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst5 (.I0(I0[5]), .I1(I1[5]), .I2(1'b0), .I3(1'b0), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst6 (.I0(I0[6]), .I1(I1[6]), .I2(1'b0), .I3(1'b0), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst7 (.I0(I0[7]), .I1(I1[7]), .I2(1'b0), .I3(1'b0), .O(inst7_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst8 (.I0(I0[8]), .I1(I1[8]), .I2(1'b0), .I3(1'b0), .O(inst8_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst9 (.I0(I0[9]), .I1(I1[9]), .I2(1'b0), .I3(1'b0), .O(inst9_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst10 (.I0(I0[10]), .I1(I1[10]), .I2(1'b0), .I3(1'b0), .O(inst10_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst11 (.I0(I0[11]), .I1(I1[11]), .I2(1'b0), .I3(1'b0), .O(inst11_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst12 (.I0(I0[12]), .I1(I1[12]), .I2(1'b0), .I3(1'b0), .O(inst12_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst13 (.I0(I0[13]), .I1(I1[13]), .I2(1'b0), .I3(1'b0), .O(inst13_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst14 (.I0(I0[14]), .I1(I1[14]), .I2(1'b0), .I3(1'b0), .O(inst14_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst15 (.I0(I0[15]), .I1(I1[15]), .I2(1'b0), .I3(1'b0), .O(inst15_O));
assign O = {inst15_O,inst14_O,inst13_O,inst12_O,inst11_O,inst10_O,inst9_O,inst8_O,inst7_O,inst6_O,inst5_O,inst4_O,inst3_O,inst2_O,inst1_O,inst0_O};
endmodule

module main (input [7:0] J1, output [7:0] J3, input  CLKIN);
wire [15:0] inst0_RDATA;
wire  inst1_O;
wire  inst2_O;
wire  inst3_O;
wire  inst4_O;
wire  inst5_O;
wire  inst6_O;
wire  inst7_O;
wire  inst8_Q;
wire  inst9_O;
wire  inst10_O;
wire [7:0] inst11_O;
wire [7:0] inst12_O;
wire  inst12_COUT;
wire [7:0] inst13_O;
wire [7:0] inst14_O;
wire [7:0] inst15_O;
wire [7:0] inst16_O;
wire [7:0] inst17_O;
wire [7:0] inst18_O;
wire [7:0] inst19_O;
wire [7:0] inst20_O;
wire [7:0] inst21_O;
wire [7:0] inst22_O;
wire [7:0] inst23_O;
wire [7:0] inst24_O;
wire [7:0] inst25_O;
wire [7:0] inst26_O;
wire [7:0] inst27_O;
wire [7:0] inst28_O;
wire [7:0] inst29_O;
wire [7:0] inst30_O;
wire [7:0] inst31_O;
wire [15:0] inst32_O;
wire [15:0] inst33_O;
wire [7:0] inst34_O;
wire [7:0] inst35_O;
wire [7:0] inst36_O;
wire [7:0] inst37_O;
wire [7:0] inst38_O;
wire [7:0] inst39_O;
wire [7:0] inst40_O;
wire [7:0] inst41_O;
wire [7:0] inst42_O;
wire [7:0] inst43_O;
wire [7:0] inst44_O;
wire [7:0] inst45_O;
wire [7:0] inst46_O;
wire [7:0] inst47_O;
wire [7:0] inst48_O;
wire [7:0] inst49_O;
wire [7:0] inst50_O;
wire [7:0] inst51_O;
wire [7:0] inst52_O;
wire [7:0] inst53_O;
wire [7:0] inst54_O;
wire [7:0] inst55_O;
wire [7:0] inst56_O;
wire [7:0] inst57_O;
wire [7:0] inst58_O;
wire [7:0] inst59_O;
wire [7:0] inst60_O;
wire [7:0] inst61_O;
wire [7:0] inst62_O;
wire [7:0] inst63_O;
wire  inst64_O;
wire [7:0] inst65_O;
wire  inst66_O;
SB_RAM40_4K #(.INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_0(256'h0000000000000000000000000000000000000000000000000000CF00B0008055),
.INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
.READ_MODE(0),
.INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
.INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000),
.WRITE_MODE(0),
.INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000)) inst0 (.RDATA(inst0_RDATA), .RADDR({1'b0,1'b0,1'b0,inst11_O[7],inst11_O[6],inst11_O[5],inst11_O[4],inst11_O[3],inst11_O[2],inst11_O[1],inst11_O[0]}), .RCLK(CLKIN), .RCLKE(1'b1), .RE(1'b1), .WCLK(CLKIN), .WCLKE(1'b0), .WE(1'b0), .WADDR({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .MASK({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}), .WDATA({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}));
SB_LUT4 #(.LUT_INIT(16'h0001)) inst1 (.I0(inst0_RDATA[14]), .I1(inst0_RDATA[15]), .I2(1'b0), .I3(1'b0), .O(inst1_O));
SB_LUT4 #(.LUT_INIT(16'h0002)) inst2 (.I0(inst0_RDATA[14]), .I1(inst0_RDATA[15]), .I2(1'b0), .I3(1'b0), .O(inst2_O));
SB_LUT4 #(.LUT_INIT(16'h0003)) inst3 (.I0(inst0_RDATA[14]), .I1(inst0_RDATA[15]), .I2(1'b0), .I3(1'b0), .O(inst3_O));
SB_LUT4 #(.LUT_INIT(16'h0100)) inst4 (.I0(inst0_RDATA[12]), .I1(inst0_RDATA[13]), .I2(inst0_RDATA[14]), .I3(inst0_RDATA[15]), .O(inst4_O));
SB_LUT4 #(.LUT_INIT(16'h0400)) inst5 (.I0(inst0_RDATA[12]), .I1(inst0_RDATA[13]), .I2(inst0_RDATA[14]), .I3(inst0_RDATA[15]), .O(inst5_O));
SB_LUT4 #(.LUT_INIT(16'h0800)) inst6 (.I0(inst0_RDATA[12]), .I1(inst0_RDATA[13]), .I2(inst0_RDATA[14]), .I3(inst0_RDATA[15]), .O(inst6_O));
SB_LUT4 #(.LUT_INIT(16'h1000)) inst7 (.I0(inst0_RDATA[12]), .I1(inst0_RDATA[13]), .I2(inst0_RDATA[14]), .I3(inst0_RDATA[15]), .O(inst7_O));
SB_DFF inst8 (.C(CLKIN), .D(inst9_O), .Q(inst8_Q));
SB_LUT4 #(.LUT_INIT(16'h6666)) inst9 (.I0(inst8_Q), .I1(1'b1), .I2(1'b0), .I3(1'b0), .O(inst9_O));
SB_LUT4 #(.LUT_INIT(16'hFE00)) inst10 (.I0(inst3_O), .I1(inst4_O), .I2(inst5_O), .I3(inst8_Q), .O(inst10_O));
Register8CE inst11 (.I(inst13_O), .O(inst11_O), .CLK(CLKIN), .CE(inst8_Q));
Add8 inst12 (.I0(inst11_O), .I1({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b1}), .O(inst12_O), .COUT(inst12_COUT));
Mux2x8 inst13 (.I0(inst12_O), .I1({inst0_RDATA[7],inst0_RDATA[6],inst0_RDATA[5],inst0_RDATA[4],inst0_RDATA[3],inst0_RDATA[2],inst0_RDATA[1],inst0_RDATA[0]}), .S(inst7_O), .O(inst13_O));
Mux2x8 inst14 (.I0({inst0_RDATA[7],inst0_RDATA[6],inst0_RDATA[5],inst0_RDATA[4],inst0_RDATA[3],inst0_RDATA[2],inst0_RDATA[1],inst0_RDATA[0]}), .I1(J1), .S(inst5_O), .O(inst14_O));
Mux2x8 inst15 (.I0(inst63_O), .I1(inst14_O), .S(inst64_O), .O(inst15_O));
Register8CE inst16 (.I(inst15_O), .O(inst16_O), .CLK(CLKIN), .CE(inst33_O[0]));
Register8CE inst17 (.I(inst15_O), .O(inst17_O), .CLK(CLKIN), .CE(inst33_O[1]));
Register8CE inst18 (.I(inst15_O), .O(inst18_O), .CLK(CLKIN), .CE(inst33_O[2]));
Register8CE inst19 (.I(inst15_O), .O(inst19_O), .CLK(CLKIN), .CE(inst33_O[3]));
Register8CE inst20 (.I(inst15_O), .O(inst20_O), .CLK(CLKIN), .CE(inst33_O[4]));
Register8CE inst21 (.I(inst15_O), .O(inst21_O), .CLK(CLKIN), .CE(inst33_O[5]));
Register8CE inst22 (.I(inst15_O), .O(inst22_O), .CLK(CLKIN), .CE(inst33_O[6]));
Register8CE inst23 (.I(inst15_O), .O(inst23_O), .CLK(CLKIN), .CE(inst33_O[7]));
Register8CE inst24 (.I(inst15_O), .O(inst24_O), .CLK(CLKIN), .CE(inst33_O[8]));
Register8CE inst25 (.I(inst15_O), .O(inst25_O), .CLK(CLKIN), .CE(inst33_O[9]));
Register8CE inst26 (.I(inst15_O), .O(inst26_O), .CLK(CLKIN), .CE(inst33_O[10]));
Register8CE inst27 (.I(inst15_O), .O(inst27_O), .CLK(CLKIN), .CE(inst33_O[11]));
Register8CE inst28 (.I(inst15_O), .O(inst28_O), .CLK(CLKIN), .CE(inst33_O[12]));
Register8CE inst29 (.I(inst15_O), .O(inst29_O), .CLK(CLKIN), .CE(inst33_O[13]));
Register8CE inst30 (.I(inst15_O), .O(inst30_O), .CLK(CLKIN), .CE(inst33_O[14]));
Register8CE inst31 (.I(inst15_O), .O(inst31_O), .CLK(CLKIN), .CE(inst33_O[15]));
Decoder4 inst32 (.I({inst0_RDATA[11],inst0_RDATA[10],inst0_RDATA[9],inst0_RDATA[8]}), .O(inst32_O));
And2x16 inst33 (.I0(inst32_O), .I1({inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O,inst10_O}), .O(inst33_O));
Mux2x8 inst34 (.I0(inst16_O), .I1(inst17_O), .S(inst0_RDATA[8]), .O(inst34_O));
Mux2x8 inst35 (.I0(inst18_O), .I1(inst19_O), .S(inst0_RDATA[8]), .O(inst35_O));
Mux2x8 inst36 (.I0(inst20_O), .I1(inst21_O), .S(inst0_RDATA[8]), .O(inst36_O));
Mux2x8 inst37 (.I0(inst22_O), .I1(inst23_O), .S(inst0_RDATA[8]), .O(inst37_O));
Mux2x8 inst38 (.I0(inst24_O), .I1(inst25_O), .S(inst0_RDATA[8]), .O(inst38_O));
Mux2x8 inst39 (.I0(inst26_O), .I1(inst27_O), .S(inst0_RDATA[8]), .O(inst39_O));
Mux2x8 inst40 (.I0(inst28_O), .I1(inst29_O), .S(inst0_RDATA[8]), .O(inst40_O));
Mux2x8 inst41 (.I0(inst30_O), .I1(inst31_O), .S(inst0_RDATA[8]), .O(inst41_O));
Mux2x8 inst42 (.I0(inst34_O), .I1(inst35_O), .S(inst0_RDATA[9]), .O(inst42_O));
Mux2x8 inst43 (.I0(inst36_O), .I1(inst37_O), .S(inst0_RDATA[9]), .O(inst43_O));
Mux2x8 inst44 (.I0(inst38_O), .I1(inst39_O), .S(inst0_RDATA[9]), .O(inst44_O));
Mux2x8 inst45 (.I0(inst40_O), .I1(inst41_O), .S(inst0_RDATA[9]), .O(inst45_O));
Mux2x8 inst46 (.I0(inst42_O), .I1(inst43_O), .S(inst0_RDATA[10]), .O(inst46_O));
Mux2x8 inst47 (.I0(inst44_O), .I1(inst45_O), .S(inst0_RDATA[10]), .O(inst47_O));
Mux2x8 inst48 (.I0(inst46_O), .I1(inst47_O), .S(inst0_RDATA[11]), .O(inst48_O));
Mux2x8 inst49 (.I0(inst16_O), .I1(inst17_O), .S(inst0_RDATA[4]), .O(inst49_O));
Mux2x8 inst50 (.I0(inst18_O), .I1(inst19_O), .S(inst0_RDATA[4]), .O(inst50_O));
Mux2x8 inst51 (.I0(inst20_O), .I1(inst21_O), .S(inst0_RDATA[4]), .O(inst51_O));
Mux2x8 inst52 (.I0(inst22_O), .I1(inst23_O), .S(inst0_RDATA[4]), .O(inst52_O));
Mux2x8 inst53 (.I0(inst24_O), .I1(inst25_O), .S(inst0_RDATA[4]), .O(inst53_O));
Mux2x8 inst54 (.I0(inst26_O), .I1(inst27_O), .S(inst0_RDATA[4]), .O(inst54_O));
Mux2x8 inst55 (.I0(inst28_O), .I1(inst29_O), .S(inst0_RDATA[4]), .O(inst55_O));
Mux2x8 inst56 (.I0(inst30_O), .I1(inst31_O), .S(inst0_RDATA[4]), .O(inst56_O));
Mux2x8 inst57 (.I0(inst49_O), .I1(inst50_O), .S(inst0_RDATA[5]), .O(inst57_O));
Mux2x8 inst58 (.I0(inst51_O), .I1(inst52_O), .S(inst0_RDATA[5]), .O(inst58_O));
Mux2x8 inst59 (.I0(inst53_O), .I1(inst54_O), .S(inst0_RDATA[5]), .O(inst59_O));
Mux2x8 inst60 (.I0(inst55_O), .I1(inst56_O), .S(inst0_RDATA[5]), .O(inst60_O));
Mux2x8 inst61 (.I0(inst57_O), .I1(inst58_O), .S(inst0_RDATA[6]), .O(inst61_O));
Mux2x8 inst62 (.I0(inst59_O), .I1(inst60_O), .S(inst0_RDATA[6]), .O(inst62_O));
Mux2x8 inst63 (.I0(inst61_O), .I1(inst62_O), .S(inst0_RDATA[7]), .O(inst63_O));
SB_LUT4 #(.LUT_INIT(16'hEEEE)) inst64 (.I0(inst5_O), .I1(inst4_O), .I2(1'b0), .I3(1'b0), .O(inst64_O));
Register8CE inst65 (.I(inst48_O), .O(inst65_O), .CLK(CLKIN), .CE(inst66_O));
SB_LUT4 #(.LUT_INIT(16'h8888)) inst66 (.I0(inst6_O), .I1(inst8_Q), .I2(1'b0), .I3(1'b0), .O(inst66_O));
assign J3 = inst65_O;
endmodule

